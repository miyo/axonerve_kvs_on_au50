`define OPT_DATA_W
//`define HBM_PRBS_ADDR_WIDTH_28
//`define HBM_PRBS_ADDR_WIDTH_27
`define HBM_PRBS_ADDR_WIDTH_23
`define P_HBM_SCH_EN_0
`define P_HBM_SCH_EN_1
